entity HALF_ADDER is
  port(
    A, B: in bit;
    SUM, CARRY: out bit);
end entity HALF_ADDER;
