architecture RTL of HALF_ADDER is
begin
  SUM <= A xor B;
  CARRY <= A and B;
end architecture RTL;
